`ifndef RKV_AHBRAM_PKG_SV
`define RKV_AHBRAM_PKG_SV

package rkv_ahbram_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  import lvc_ahb_pkg::*;

endpackage



`endif // RKV_AHBRAM_PKG_SV
