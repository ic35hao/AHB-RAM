
module rkv_ahbram_tb;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  import rkv_ahbram_pkg::*;

  ahb_blockram_32 dut();

  initial begin
    //run_test();
  end


endmodule
