`ifndef RKV_AHBRAM_SEQ_LIB_SVH
`define RKV_AHBRAM_SEQ_LIB_SVH

`include "rkv_ahbram_element_sequences.svh"
`include "rkv_ahbram_base_virtual_sequence.sv"
`include "rkv_ahbram_smoke_virt_seq.sv"


`endif
