`ifndef RKV_AHBRAM_IF_SV
`define RKV_AHBRAM_IF_SV

interface rkv_ahbram_if;
  logic clk;
  logic rstn;

endinterface


`endif // RKV_AHBRAM_IF_SV

